`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: BIT
// Engineer: ZHC
// 
// Create Date: 2020/09/10 09:56:56
// Design Name: 
// Module Name: ALU
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////

module ALU(
	input [11:0] alu_op,
	input [31:0] alu_src1,
	input [31:0] alu_src2,
	output [31:0] alu_result
	);
	//�������в�����
	wire op_add;	//�ӷ�
	wire op_sub;	//����
	wire op_slt;	//�з������Ƚϣ�С����1
	wire op_sltu;	//�޷������Ƚϣ�С����1
	wire op_and;	//��λ��
	wire op_nor;	//��λ���
	wire op_or;		//��λ��
	wire op_xor;	//��λ���
	wire op_sll;	//�߼�����
	wire op_srl;	//�߼�����
	wire op_sra;	//��������
	wire op_lui;	//���������ڸ߰벿��

	//Ϊ���в�������ֵ
	assign op_add 	= alu_op[ 0];
	assign op_sub 	= alu_op[ 1];
	assign op_slt 	= alu_op[ 2];
	assign op_sltu 	= alu_op[ 3];
	assign op_and 	= alu_op[ 4];
	assign op_nor 	= alu_op[ 5];
	assign op_or 	= alu_op[ 6];
	assign op_xor 	= alu_op[ 7];
	assign op_sll 	= alu_op[ 8];
	assign op_srl 	= alu_op[ 9];
	assign op_sra 	= alu_op[10];
	assign op_lui 	= alu_op[11];

	//�������н��
	wire [31:0] add_sub_result;
	wire [31:0] slt_result;
	wire [31:0] sltu_result;
	wire [31:0] and_result;
	wire [31:0] nor_result;
	wire [31:0] or_result;
	wire [31:0] xor_result;
	wire [31:0] lui_result;
	wire [31:0] sll_result;
	wire [31:0] sr64_result;
	wire [31:0] sr_result;

	//�����м����
	wire [31:0] adder_a;
	wire [31:0] adder_b;
	wire 		adder_cin;
	wire [31:0] adder_result;
	wire 		adder_cout;

	/*ʵ�ּӼ���*/
	assign adder_a = alu_src1;
	assign adder_b = (op_sub | op_slt | op_sltu) ? ~alu_src2 : alu_src2; 
	//����Ǽ�������ȡ�����ټ�1�õ�����
	assign adder_cin = (op_sub | op_slt | op_sltu) ? 1'b1 : 1'b0;
	assign {adder_cout, adder_result} = adder_a + adder_b + adder_cin;
	assign add_sub_result = adder_result;

	/*ʵ���з������޷������ıȽ�*/
	assign slt_result[31:1] = 31'b0;
	//����������һ��һ����������������ͬ�Ž��Ϊ����
	assign slt_result[0] = (alu_src1[31] & ~alu_src2[31])
							| ((~alu_src1[31] ^ alu_src2[31]) & adder_result[31]);
	//�޷�������ӣ��޽�λ��˵��С��
	assign sltu_result[31:1] = 31'b0;
	assign sltu_result[0] = ~adder_cout;

	/*ʵ��λ����*/
	assign and_result = alu_src1 & alu_src2;
	assign or_result = alu_src1 | alu_src2;
	assign nor_result = ~or_result;
	assign xor_result = alu_src1 ^ alu_src2;

	assign lui_result = {alu_src2[15:0], 16'b0};

	/*ʵ����������*/
	assign sll_result = alu_src2 << alu_src1[4:0];
	//�����sra�����Ʋ������λ�������srl�����Ʋ���0
	assign sr64_result = {{32{op_sra & alu_src2[31]}}, alu_src2[31:0]} >> alu_src1[4:0];
	assign sr_result = sr64_result[31:0];

	//���Ķ�·ѡ����
	assign alu_result = ({32{op_add | op_sub}} & add_sub_result)
				  	  | ({32{op_slt}} & slt_result)
				  	  | ({32{op_sltu}} & sltu_result)
				  	  | ({32{op_and}} & and_result)
				  	  | ({32{op_nor}} & nor_result)
				  	  | ({32{op_or}} & or_result)
				  	  | ({32{op_xor}} & xor_result)
				  	  | ({32{op_lui}} & lui_result)
				  	  | ({32{op_sll}} & sll_result)
				  	  | ({32{op_sra | op_srl}} & sr_result);
endmodule
